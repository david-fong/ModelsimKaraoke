`define CHAR_H 9
`define CHAR_W 6
`define CHAR_N 600
`define ADDR_W 12