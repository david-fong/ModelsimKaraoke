`define CHAR_H 9
`define CHAR_W 6
`define LINE_N 22
`define CPSBLN 24
`define CHAR_W 6
`define ADDR_W 16
