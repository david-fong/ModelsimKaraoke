`define CHAR_H 9
`define CHAR_W 6
`define LINE_N 49
`define CPSBLN 21
`define CHAR_W 6
`define ADDR_W 32
